//(c) Alina Ivanova, alina.al.ivanova@gmail.com
//----------------------------------------------------------------------------- 
package package_settings;
//-----------------------------------------------------------------------------
// Parameter Declaration(s)
//-----------------------------------------------------------------------------
	parameter SIZE_MAX_WINDOW                 = 64;
	parameter SIZE_WINDOW                     = 8;
	parameter SIZE_DATA                       = 16;
//-----------------------------------------------------------------------------
endpackage: package_settings
