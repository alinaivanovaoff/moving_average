//-----------------------------------------------------------------------------
// Title       : package_settings (parameters)
//-----------------------------------------------------------------------------
// File        : package_settings.sv
// Company     : My company
// Created     : 11/03/2014
// Created by  : Alina Ivanova
//-----------------------------------------------------------------------------
// Description : settings package
//-----------------------------------------------------------------------------
// Revision    : 1.0
//-----------------------------------------------------------------------------
// Copyright (c) 2014 My company
// This work may not be copied, modified, re-published, uploaded, executed, or
// distributed in any way, in any medium, whether in whole or in part, without
// prior written permission from My Company.
//-----------------------------------------------------------------------------
//-----------------------------------------------------------------------------
package package_settings;
//-----------------------------------------------------------------------------
// Parameter Declaration(s)
//-----------------------------------------------------------------------------
	parameter SIZE_MAX_WINDOW                 = 64;
	parameter SIZE_WINDOW                     = 8;
	parameter SIZE_DATA                       = 16;
//-----------------------------------------------------------------------------
//-----------------------------------------------------------------------------
endpackage
